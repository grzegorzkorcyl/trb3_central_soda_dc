-------------------------------------
-- Defines the dataPath width
--
-------------------------------------
package mypackage is
   constant XBITS :INTEGER := 32; 
   constant YBITS :INTEGER := 32;
   constant GRAIN :INTEGER := 2; --Allways in 2!!!!
   constant DEPTH :INTEGER := 1; --Every how much steps register
end mypackage;
