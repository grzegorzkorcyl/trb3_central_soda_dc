----------------------------------------------------------------------------------
-- Company:       KVI/RUG/Groningen University
-- Engineer:      Peter Schakel
-- Create Date:   12-07-2013
-- Module Name:   DC_module_TRB3
-- Description:   Multiplexer module for TRB3
-- Modifications:
--   30-07-2014   Timestamp from FEE is now composed by 16 bits superburstnumber and timestamp counter within superburst
--   29-08-2014   ADCCLOCKFREQUENCY added: SODA clock at 80MHz 
--   27-01-2015   SCI interface removed
--   28-01-2015   Histogram removed
--   26-02-2015   added signal no_packet_limit for unlimited data output
--   21-05-2015   Moved serdes/gtx part to top-level
--   21-05-2015   Additional clock synchronization
--   15-09-2015   Sorting waveform multiplexer instead of unsorted
--   02-10-2015   Sorting hit multiplexer input now with hit-data members instead of 36-bits data
----------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.all ;
USE ieee.std_logic_arith.all ;
USE work.panda_package.all;

----------------------------------------------------------------------------------
-- DC_module_TRB3
-- Module to describe the behavioral of the Panda Data collector multiplexer.
-- Soda signals are generated by a SODA generator.
-- Slow control is done by TRBnet.
--    
-- Connection to the Front End Electronics fibers is implemented with synchronized serdes fiber link:
-- From MUX to FEE the clock is phase aligned for SODA signals. Asynchronous data is used for slow control.
-- From FEE to MUX the clock is not phase aligned. The connection is used for pulse data and slow control.
-- Pulse data from the FEE fiber data is available in packets of 4*36-bits words.
-- The pulse data from the fibres are combined to one stream. The pulse-data is sorted on the timestamp and the time-fraction.
-- The pileup waveform data from the fibres are also combined to one stream. This is not sorted.
-- The resulting streams with pulse data and with pileup waveforms are combined into 64-bit data according to Panda data format.
--
-- Adresses from slowcontrol module, see work.panda_package for constants:
--     ADDRESS_MUX_SODA_CONTROL :
--         only write: settings for the SODA : 
--         bit0 : enable SODA packets
--         bit1 : reset timestamp counters
--         bit2 : Enable data taking 
--         bit3 : Disable data taking
--         bit4 : Enable 64-bit output data
--         bit5 : Enable Pileup Waveform sending
--         bit6 : Select source for multiplexer status (ADDRESS_MUX_MULTIPLEXER_STATUS): 0=pulse, 1=waveform
--
--     ADDRESS_MUX_EXTRACTWAVE
--         request: start extracting waveform of 1 pileup pulse:
--         bit 15..0 : selected adcnumber (if bit 16 is set)
--         bit 16 : select 1 adc, otherwise take first data arriving
--         bit 17 : select 1 low/high combination instead of 1 adc channel
--         The reply will be (after a waveform has been measured) :
--         32-bits word0  : bits(31..24)=0xD0, bits23..0=ADDRESS_MUX_EXTRACTWAVE
--         32-bits word1  : bits(31..0)=timestamp of maximum value in waveform
--         32-bits word2  : bits(31)=0, bits(30..0)=SuperBurst number
--         32-bits word3  : bits(31..24) = statusbyte, bits(23..16) = 00, bits(15..0) = adcnumber 
--         32-bits word4..n: bit(31)=0, bits(30..16)=adc sample, bit(15)=0, bits(14..0)=next adc sample
--         32-bits last word (1sample): bits(31)=1, bits(30..16)=last adc sample, bit(15)=0, bits(14..0)=0
--         32-bits last word (2samples): bits(31)=0, bits(30..16)=adc sample, bit15=1, bits(14..0)=last adc sample
--         32-bits last word (error): bits(31)=1, bits(30..16)=don't care, bit15=1, bits(14..0)=don't care
--
--     ADDRESS_MUX_EXTRACTDATA
--         request: start extracting data of 1 pulse:
--         bit 15..0 : selected adcnumber
--         bit 16 : select 1 adc, otherwise take first data arriving
--         bit 17 : select 1 low/high combination instead of 1 adc channel
--         The reply will be :
--         32-bits word0  : bits(31..24=0xD0, bits23..0=ADDRESS_MUX_EXTRACTDATA
--         32-bits word1  : bits(31..24)=statusbyte, bits(23..16)=0, bits(15..0)=adcnumber
--         32-bits word2  : bits(31..24)=0xD0, bits(23..0)=ADDRESS_MUX_EXTRACTDATA+1
--         32-bits word3  : bits(31..24)=timefraction, bits(15..0)=energy
--         32-bits word4  : bits(31..24)=0xD0, bits(23..0)= ADDRESS_MUX_EXTRACTDATA+2
--         32-bits word5  : bits(31..0)= timestamp(47..16) with bits 47..32 set to 0
--         32-bits word6  : bits(31..24)=0xD0, bits23..0= ADDRESS_MUX_EXTRACTDATA+3
--         32-bits word7  : bits(31..16)=0, bits(15..0)=timestamp(15..0)
--
--     ADDRESS_MUX_SYSMON
--         write to FPGA system monitor
--         bit 31 : slect read/write, write='0', read='1'
--         bit 30 : reset/reconfigure FPGA system monitor
--         bit 22..16 : 7-bits address of FPGA system monitor
--         bit 15..0 : 16-bits data for FPGA system monitor
--         read from FPGA system monitor, effective address is the last address at data bits 30..16 that was written
--         bit 30..16 : 7-bits effective address of FPGA system monitor
--         bit 15..0 : data from FPGA system monitor
--
--
-- Library
--     work.panda_package :  for type declarations and constants
-- 
-- Generics:
--     NROFFIBERS : number of fiber connection of the MUX board (only 4 is possible)
--     NROFADCS : number of ADCs in each FEE
--     ADCBITS : number of analog to digital conversion bits
--     ADCCLOCKFREQUENCY : Frequency of the ADCclock in Hz, defines also the SODA clock frequency
--     MAX_DIVIDERSCALEBITS : number of scaling bits for division two largest samples
--     MAX_LUTSIZEBITS : number of bits the maximum correction Look Up Table
--     MAX_LUTSCALEBITS : number of scaling bits for the correction on the maximum (energy)
--     MUXINFIFOSIZE : size (fifo-depth bits) of the input fifo's of the multiplexer
--     TRANSFERFIFOSIZE : size (fifo-depth bits) of multiplexer transfer fifo
--     CF_FRACTIONBIT : number of valid constant fraction bits
--     TRANSITIONBUFFERBITS : number of bits for the buffer that stores data from the next superburst
--     PANDAPACKETBUFFERBITS : number of bits for the buffer to store packet for size calculation
--     ADCINDEXSHIFT : ADC channel numbers lowest bit indicates the high or low gain ADC, 0=high, 1=low
--     ENERGYSCALINGBITS : number of scaling bits for energy adjustment: energy = (original_energy * gainfactor<<scalingbits)>>scalingbits
--     COMBINEPULSESMEMSIZE : addressbits for the fifo buffer for combining hits
--     COMBINETIMEDIFFERENCE : largest time difference between hits to be combined, number of timefraction units
--     SYSTEM_ID : ID number of this Data Concentrator
-- 
-- Inputs:
--     slowcontrol_clock : clock for the slowcontrol input/output
--     packet_in_clock : clock for data from the fiber module
--     MUX_clock : clock for the multiplexer
--     packet_out_clock : clock for data from the multiplexer output
--     SODA_clock : clock for SODA signals
--     reset : reset of all components
--     BUS_READ_IN : TRBnet local bus read signal
--     BUS_WRITE_IN : TRBnet local bus write signal
--     BUS_ADDR_IN : TRBnet local bus address
--     BUS_DATA_IN : TRBnet local bus data
--     fiber_txlocked : lock signal from fiber transmitter
--     fiber_rxlocked : lock signal from fiber receiver
--     fiber_data32fifofull : fifo of fiber transmitter is full
--     fiber_data32present : fifo of fiber receiver has data available
--     fiber_data32in : 32 bits data from fiber receiver
--     fiber_rxerror : error in received data from fiber
--     superburst_number : actual superburst number received from SODA
--     superburst_update : signal for new superburst number received from SODA
--     data_out_allowed : 64-bits output data allowed to write (normally: connected fifo not full)
-- 
-- Outputs:
--     BUS_BUSY_OUT : TRBnet local bus busy signal
--     BUS_ACK_OUT : TRBnet local bus acknowledge signal
--     BUS_DATA_OUT : TRBnet local bus data
--     reset_fibers : reset fiber receiver/transmitters
--     fiber_data32write : write signal for 32bits data to fiber transmitter
--     fiber_data32out : 32bits data to fiber transmitter
--     fiber_data32read : read signal for 32bits data from fiber receiver
--     SODA_enable : enable signal for SODA receiver/transmitter
--     EnableExternalSODA : Enable external (fibre coupled) SODA instead of internal SODA generation (for debugging, not used)
--     data_out : 64-bits output data
--     data_out_write : 64-bits output data write signal
--     data_out_first : 64-bits output data first word in packet
--     data_out_last : 64-bits output data last word in packet
--     data_out_error : error occured in 64-bits output data
--     no_packet_limit : control signal for unlimited data throughput (minimum time between packets)
-- 
-- Components:
--     DC_slow_control_TRB3 : module for slow control : TRBnet local bus to Data Concentrator registers/status
--     DC_posedge_to_pulse : Makes a 1-clock pulse on rising edge from signal with different clock
--     DC_Quad_fiber_module : Handles the connection to/from the FEE, builds & entangles fiber packets (for one module for 4 fibers)
--     DC_sorting_mux : Multiplex the pulse data from all the fiber inputs to one output and sort it based on timestamp
--     DC_wavemux : Multiplex the pileup waveform data from all the fiber inputs to one output
--     DC_check_timestamp : check if the timestamps are sorted well
--     DC_extract_data : Extract pulse data from the data stream for handling by slow control
--     DC_extract_wave : Extract pileup waveform from the data stream for handling by slow control
--     DC_data_wave_to_64bit : put pulse and waveform data in packets with 64-bits wide bus
--     DC_combine_pulses : Combine pulses (=hits) from corresponding ADC channels
--     sync_bit : Synchronization for 1 bit cross clock signal
--
----------------------------------------------------------------------------------

entity DC_module_TRB3 is
	generic (
		NROFFIBERS              : natural := 4;
		NROFADCS                : natural := 16;
		ADCBITS                 : natural := 14;
		ADCCLOCKFREQUENCY       : natural := 80000000;
		MAX_DIVIDERSCALEBITS    : natural := 12;
		MAX_LUTSIZEBITS         : natural := 8;
		MAX_LUTSCALEBITS        : natural := 14;
		MUXINFIFOSIZE           : natural := 9;
		TRANSFERFIFOSIZE        : natural := 14;
		CF_FRACTIONBIT          : natural := 11;
		TRANSITIONBUFFERBITS    : natural := 7;
		PANDAPACKETBUFFERBITS   : natural := 13;
		ADCINDEXSHIFT           : natural := 1;
		ENERGYSCALINGBITS       : natural := 13;
		COMBINEPULSESMEMSIZE    : natural := 10;
		COMBINETIMEDIFFERENCE   : natural := 5000;
		SYSTEM_ID               : std_logic_vector(15 downto 0) := x"5555"		
	);
	port ( 
		slowcontrol_clock       : in std_logic;
		packet_in_clock         : in std_logic;
		MUX_clock               : in std_logic;
		packet_out_clock        : in std_logic;
		SODA_clock              : in std_logic;
		reset                   : in std_logic;

-- Slave bus
		BUS_READ_IN             : in   std_logic;
		BUS_WRITE_IN            : in   std_logic;
		BUS_BUSY_OUT            : out  std_logic;
		BUS_ACK_OUT             : out  std_logic;
		BUS_ADDR_IN             : in   std_logic_vector(1 downto 0);
		BUS_DATA_IN             : in   std_logic_vector(31 downto 0);
		BUS_DATA_OUT            : out  std_logic_vector(31 downto 0);
		
-- fiber interface signals:
		fiber_txlocked          : in std_logic_vector(0 to NROFFIBERS-1);
		fiber_rxlocked          : in std_logic_vector(0 to NROFFIBERS-1);
		reset_fibers            : out std_logic;
		fiber_data32write       : out std_logic_vector(0 to NROFFIBERS-1);
		fiber_data32out         : out array_fiber32bits_type;
		fiber_data32fifofull    : in std_logic_vector(0 to NROFFIBERS-1);
		fiber_data32read        : out std_logic_vector(0 to NROFFIBERS-1);
		fiber_data32present     : in std_logic_vector(0 to NROFFIBERS-1);
		fiber_data32in          : in array_fiber32bits_type;
		fiber_rxerror           : in std_logic_vector(0 to NROFFIBERS-1);
			
-- SODA signals
		superburst_number       : in std_logic_vector(30 downto 0);
		superburst_update       : in std_logic;
		SODA_enable             : out std_logic;
		EnableExternalSODA      : out std_logic;

-- 64 bits data output
		data_out_allowed        : in std_logic;
		data_out                : out std_logic_vector(63 downto 0);
		data_out_write          : out std_logic;
		data_out_first          : out std_logic;
		data_out_last           : out std_logic;
		data_out_error          : out std_logic;
		no_packet_limit         : out std_logic;
		
-- testpoints
		testword0               : out std_logic_vector (35 downto 0) := (others => '0');
		testword0clock          : out std_logic := '0';
		testword1               : out std_logic_vector (35 downto 0) := (others => '0');
		testword2               : out std_logic_vector (35 downto 0) := (others => '0')

		);
end DC_module_TRB3;

architecture Behavioral of DC_module_TRB3 is

component DC_slow_control_TRB3 is
	port(	
		rst                     : in std_logic;
		clk                     : in std_logic;
-- Slave bus
		BUS_READ_IN             : in   std_logic;
		BUS_WRITE_IN            : in   std_logic;
		BUS_BUSY_OUT            : out  std_logic;
		BUS_ACK_OUT             : out  std_logic;
		BUS_ADDR_IN             : in   std_logic_vector(1 downto 0);
		BUS_DATA_IN             : in   std_logic_vector(31 downto 0);
		BUS_DATA_OUT            : out  std_logic_vector(31 downto 0);

		io_data_in              : in std_logic_vector(0 to NROFFIBERS-1);
		IO_data_in_available    : in std_logic_vector(0 to NROFFIBERS-1);
		io_data_out             : out std_logic_vector(7 downto 0);
		io_write_out            : out std_logic;

		extract_data_available  : in std_logic;
		extract_wave_available  : in std_logic;

		board_status            : in array_muxregister_type;
		board_status_read       : out std_logic_vector(0 to NROFMUXREGS-1);
		board_control           : out array_muxregister_type;
		board_control_write     : out std_logic_vector(0 to NROFMUXREGS-1);
		testword0               : out std_logic_vector (35 downto 0) := (others => '0')
		);
end component;

component DC_fibermodule_interface is
	generic (
		NROFADCS                : natural := NROFADCS;
		ADCINDEXSHIFT           : natural := ADCINDEXSHIFT;
		ADCBITS                 : natural := ADCBITS;
		CF_FRACTIONBIT          : natural := CF_FRACTIONBIT;
		ENERGYSCALINGBITS       : natural := ENERGYSCALINGBITS;
		MAX_DIVIDERSCALEBITS    : natural := MAX_DIVIDERSCALEBITS;
		MAX_LUTSIZEBITS         : natural := MAX_LUTSIZEBITS;
		MAX_LUTSCALEBITS        : natural := MAX_LUTSCALEBITS
	);
	port ( 
		slowcontrol_clock       : in std_logic;
		packet_clock            : in std_logic;
		MUX_clock               : in std_logic;
		SODA_clock              : in std_logic;
		reset                   : in std_logic;
		channel                 : in std_logic_vector (3 downto 0);
		superburst_number       : in std_logic_vector(30 downto 0);
		superburst_update       : in std_logic;

-- SlowControl to/from cpu
		IO_byte                 : in std_logic_vector(7 downto 0);
		IO_write                : in std_logic;
		IO_serialdata           : out std_logic;
		IO_serialavailable      : out std_logic;
		
-- multiplexer status
		muxstat_infifo_fullness : in std_logic_vector (15 downto 0);
		muxstat_outfifo_fullness : in std_logic_vector (15 downto 0);
		timestamp_errors        : in std_logic_vector(9 downto 0);
		skipped_pulses          : in std_logic_vector(9 downto 0);
		dataerrors              : in std_logic_vector(9 downto 0);
		clearerrors             : out std_logic;
		
-- Pulse data
		channel_out             : out std_logic_vector(15 downto 0);
		statusbyte_out          : out std_logic_vector(7 downto 0);
		energy_out              : out std_logic_vector(15 downto 0);
		timefraction_out        : out std_logic_vector(11 downto 0);
		timestamp_out           : out std_logic_vector(15 downto 0);
		superburstnumber_out    : out std_logic_vector(30 downto 0);		
		pulse_data_write        : out std_logic;
		pulse_data_allowed      : in std_logic;
		pulse_data_almostfull   : in std_logic;

-- Wave data
		wave_data_out           : out std_logic_vector(35 downto 0);
		wave_data_write         : out std_logic;
		wave_data_out_allowed   : in std_logic;

-- MUX tx interface signals:
		txAsyncDataWrite        : out std_logic;
		txAsyncData             : out std_logic_vector(31 downto 0);
		txEndOfAsyncData        : out std_logic;
		txAsyncFifoFull         : in std_logic;
		txLocked                : in std_logic;

-- MUX rx interface signals:
		rxAsyncClk              : out std_logic;
		rxAsyncDataRead         : out std_logic;
		rxAsyncDataPresent      : in std_logic;
		rxAsyncData             : in std_logic_vector(31 downto 0);
		rxNotInTable            : in std_logic;
		rxLocked                : in std_logic;
		
-- Testpoints
		testword0               : out std_logic_vector (35 downto 0) := (others => '0');
		testword1               : out std_logic_vector (35 downto 0) := (others => '0')
		);
end component;

component DC_sorting_mux is
	generic(
		NROFMUXINPUTS           : natural := NROFFIBERS;
		MUXINFIFOSIZE           : natural := MUXINFIFOSIZE;
		TRANSFERFIFOSIZE        : natural := TRANSFERFIFOSIZE;
		CF_FRACTIONBIT          : natural := CF_FRACTIONBIT
	);
    port ( 
		inputclock              : in std_logic;
		MUXclock                : in std_logic; 
		outputclock             : in std_logic; 
		reset                   : in std_logic;
		channel_in              : in array_fiber16bits_type;
		statusbyte_in           : in array_fiber8bits_type;
		energy_in               : in array_fiber16bits_type;
		timefraction_in         : in array_fiber12bits_type;
		timestamp_in            : in array_fiber16bits_type;
		superburstnumber_in     : in array_fiber31bits_type;		
		data_in_write           : in std_logic_vector(0 to NROFMUXINPUTS-1);
		data_in_allowed         : out std_logic_vector(0 to NROFMUXINPUTS-1);
		data_in_almostfull      : out std_logic_vector(0 to NROFMUXINPUTS-1);
		fiber_index_out         : out std_logic_vector(3 downto 0);
		channel_out             : out std_logic_vector(15 downto 0);
		statusbyte_out          : out std_logic_vector(7 downto 0);
		energy_out              : out std_logic_vector(15 downto 0);
		timefraction_out        : out std_logic_vector(11 downto 0);
		timestamp_out           : out std_logic_vector(15 downto 0);
		superburstnumber_out    : out std_logic_vector(30 downto 0);		
		data_out_read           : in std_logic;
		data_out_available      : out std_logic;
		infifo_fullness         : out array_fiber16bits_type;
		outfifo_fullness        : out std_logic_vector(15 downto 0);
		error                   : out std_logic;
		testword0               : out std_logic_vector(35 downto 0) := (others => '0');
		testword1               : out std_logic_vector(35 downto 0) := (others => '0'));
end component;

component DC_combine_pulses is
	generic (
		NROFFIBERS              : natural := NROFFIBERS;
		NROFADCS                : natural := NROFADCS;
		ADCINDEXSHIFT           : natural := ADCINDEXSHIFT;
		COMBINEPULSESMEMSIZE    : natural := COMBINEPULSESMEMSIZE;
		COMBINETIMEDIFFERENCE   : natural := COMBINETIMEDIFFERENCE;
		CF_FRACTIONBIT          : natural := CF_FRACTIONBIT
		);
	port ( 
		clock                   : in std_logic;
		reset                   : in std_logic;
		combine_pulse           : in std_logic_vector((NROFFIBERS*NROFADCS)/(2*(ADCINDEXSHIFT+1))-1 downto 0);
		fiber_index_in          : in std_logic_vector(3 downto 0);
		channel_in              : in std_logic_vector(15 downto 0);
		statusbyte_in           : in std_logic_vector(7 downto 0);
		energy_in               : in std_logic_vector(15 downto 0);
		timefraction_in         : in std_logic_vector(11 downto 0);
		timestamp_in            : in std_logic_vector(15 downto 0);
		superburstnumber_in     : in std_logic_vector(30 downto 0);
		data_in_read            : out std_logic;
		data_in_available       : in std_logic;

		channel_out             : out std_logic_vector(15 downto 0);
		statusbyte_out          : out std_logic_vector(7 downto 0);
		energy_out              : out std_logic_vector(15 downto 0);
		timefraction_out        : out std_logic_vector(11 downto 0);
		timestamp_out           : out std_logic_vector(15 downto 0);
		superburstnumber_out    : out std_logic_vector(30 downto 0);
		data_out_read           : in std_logic;
		data_out_available      : out std_logic
	);
end component;

component DC_wavemux is
	generic(
		NROFMUXINPUTS           : natural := NROFFIBERS
	);
    Port ( 
		inputclock              : in std_logic;
		MUXclock                : in std_logic; 
		outputclock             : in std_logic; 
		reset                   : in std_logic;
		data_in                 : in array_fiber36bits_type;
		data_in_write           : in std_logic_vector(0 to NROFMUXINPUTS-1);
		data_in_wave_allowed    : out std_logic_vector(0 to NROFMUXINPUTS-1);
		data_out                : out std_logic_vector(35 downto 0);
		data_out_read           : in std_logic;
		data_out_available      : out std_logic;
		infifo_fullness         : out array_fiber16bits_type;
		outfifo_fullness        : out std_logic_vector(15 downto 0);
		testword0               : out std_logic_vector(35 downto 0) := (others => '0');
		testword1               : out std_logic_vector(35 downto 0) := (others => '0');
		error                   : out std_logic);
end component;

component DC_sorting_wavemux is
	generic(
		NROFMUXINPUTS           : natural := NROFFIBERS
	);
    Port ( 
		inputclock              : in std_logic;
		MUXclock                : in std_logic; 
		outputclock             : in std_logic; 
		reset                   : in std_logic;
		data_in                 : in array_fiber36bits_type;
		data_in_write           : in std_logic_vector(0 to NROFMUXINPUTS-1);
		data_in_wave_allowed    : out std_logic_vector(0 to NROFMUXINPUTS-1);
		data_out                : out std_logic_vector(35 downto 0);
		data_out_read           : in std_logic;
		data_out_available      : out std_logic;
		data_out_inpipe         : out std_logic;
		infifo_fullness         : out array_fiber16bits_type;
		outfifo_fullness        : out std_logic_vector(15 downto 0);
		error                   : out std_logic;
		testword0               : out std_logic_vector(35 downto 0);
		testword1               : out std_logic_vector(35 downto 0)
);
end component;

component DC_check_timestamp is
	port ( 
		clock                   : in std_logic;
		reset                   : in std_logic;
		clear                   : in std_logic;
		channel                 : in std_logic_vector(15 downto 0);
		statusbyte              : in std_logic_vector(7 downto 0);
		energy                  : in std_logic_vector(15 downto 0);
		timefraction            : in std_logic_vector(11 downto 0);
		timestamp               : in std_logic_vector(15 downto 0);
		superburstnumber        : in std_logic_vector(30 downto 0);		
		pulse_data_write        : in std_logic;
		multiplexer_error       : in std_logic;
		timestamp_errors        : out std_logic_vector(9 downto 0);	
		skipped_pulses          : out std_logic_vector(9 downto 0);
		dataerrors              : out std_logic_vector(9 downto 0)
		);
end component;

component DC_posedge_to_pulse is
	port (
		clock_in                : in  std_logic;
		clock_out               : in  std_logic;
		en_clk                  : in  std_logic;
		signal_in               : in  std_logic;
		pulse                   : out std_logic);
end component;

component DC_data_wave_to_64bit is
	generic (
		TRANSITIONBUFFERBITS : natural := TRANSITIONBUFFERBITS;
		PANDAPACKETBUFFERBITS : natural := PANDAPACKETBUFFERBITS;
		SYSTEM_ID               : std_logic_vector(15 downto 0) := SYSTEM_ID
	);
    Port ( 
		clock                   : in std_logic;
		reset                   : in std_logic;
		latestsuperburstnumber  : in std_logic_vector(30 downto 0);
		channel                 : in std_logic_vector(15 downto 0);
		statusbyte              : in std_logic_vector(7 downto 0);
		energy                  : in std_logic_vector(15 downto 0);
		timefraction            : in std_logic_vector(11 downto 0);
		timestamp               : in std_logic_vector(15 downto 0);
		superburstnumber        : in std_logic_vector(30 downto 0);		
		data_in_available       : in std_logic;
		data_in_read            : out std_logic;
		wave_in                 : in std_logic_vector(35 downto 0);
		wave_in_available       : in std_logic;
		wave_in_read            : out std_logic;
		data_out_allowed        : in std_logic;
		data_out                : out std_logic_vector(63 downto 0);
		data_out_write          : out std_logic;
		data_out_first          : out std_logic;
		data_out_last           : out std_logic;
		error                   : out std_logic;
		testword0               : out std_logic_vector(35 downto 0) := (others => '0');
		testword1               : out std_logic_vector(35 downto 0) := (others => '0')
		);
end component;

component DC_extract_data is
	port ( 
		write_clock             : in std_logic;
		read_clock              : in std_logic;
		reset                   : in std_logic;
		start                   : in std_logic;
		make_selection          : in std_logic;
		dualgain                : in std_logic;
		adcnumber               : in std_logic_vector(15 downto 0);		
		channel                 : in std_logic_vector(15 downto 0);
		statusbyte              : in std_logic_vector(7 downto 0);
		energy                  : in std_logic_vector(15 downto 0);
		timefraction            : in std_logic_vector(11 downto 0);
		timestamp               : in std_logic_vector(15 downto 0);
		superburstnumber        : in std_logic_vector(30 downto 0);		
		pulse_data_write        : in std_logic;
		ready                   : out std_logic;
		pulse_data_select       : in std_logic_vector(1 downto 0);
		pulse_data_out          : out std_logic_vector(31 downto 0);
		testword0               : out std_logic_vector(35 downto 0) := (others => '0')
		);
end component;

component DC_extract_wave is
	port ( 
		write_clock             : in std_logic;
		read_clock              : in std_logic;
		reset                   : in std_logic;
		start                   : in std_logic;
		make_selection          : in std_logic;
		dualgain                : in std_logic;
		adcnumber               : in std_logic_vector(15 downto 0);		
		wave_data_in            : in std_logic_vector(35 downto 0);
		wave_data_in_write      : in std_logic;
		ready                   : out std_logic;
		wave_data_out           : out std_logic_vector(31 downto 0);
		wave_data_out_read      : in std_logic;
		testword0               : out std_logic_vector(35 downto 0) := (others => '0')
		);
end component;

component DC_checkwave is
    Port ( 
		clock                   : in std_logic;
		reset                   : in std_logic;
		wave_in                 : in std_logic_vector(35 downto 0);
		wave_in_write           : in std_logic;
		error                   : out std_logic
	);    
end component;
constant DEBUG_SLOWCONTROL           : boolean := false;
constant ones                        : std_logic_vector(31 downto 0) := (others => '1');
signal reset_slowcontrolclock_S      : std_logic;
signal reset_packet_in_clock_S       : std_logic;
signal reset_packet_out_clock_S      : std_logic;
signal reset_SODAclock_S             : std_logic;
signal reset_fibers0_S               : std_logic;

signal EnableOutputFibre_S           : std_logic;
signal EnableOutputFibre0_S          : std_logic;
signal EnableWaveformSending_S       : std_logic;
signal SODA_TimeTagValid_S           : std_logic;

signal superburst_number_S           : std_logic_vector(30 downto 0);
signal superburst_update_S           : std_logic;

signal pulse_data_array_S            : array_fiber36bits_type := (others => (others => '0'));             
signal pulse_data_array_channel_S    : array_fiber16bits_type;
signal pulse_data_array_statusbyte_S : array_fiber8bits_type;
signal pulse_data_array_energy_S     : array_fiber16bits_type;
signal pulse_data_array_timefraction_S: array_fiber12bits_type;
signal pulse_data_array_timestamp_S  : array_fiber16bits_type;
signal pulse_data_array_superburstnumber_S: array_fiber31bits_type;		
signal pulse_data_array_write_S      : std_logic_vector (0 to NROFFIBERS-1) := (others => '0');
signal pulse_data_array_allowed_S    : std_logic_vector (0 to NROFFIBERS-1);
signal pulse_data_array_almostfull_S : std_logic_vector (0 to NROFFIBERS-1);

signal wave_data_array_S             : array_fiber36bits_type := (others => (others => '0'));                 
signal wave_data_array_write_S       : std_logic_vector (0 to NROFFIBERS-1) := (others => '0');
signal wave_data_array_allowed_S     : std_logic_vector (0 to NROFFIBERS-1);

signal wave_data_available_S         : std_logic;
signal wave_data_read_S              : std_logic;
signal wave_data_read0_S             : std_logic;
signal wave_data_S                   : std_logic_vector (35 downto 0);
signal wave_data_in_write_S          : std_logic;
--signal wave_data_read0_S             : std_logic;
		
signal fiber_index_S                 : std_logic_vector(3 downto 0);
signal mux_channel_S                 : std_logic_vector(15 downto 0);
signal mux_statusbyte_S              : std_logic_vector(7 downto 0);
signal mux_energy_S                  : std_logic_vector(15 downto 0);
signal mux_timefraction_S            : std_logic_vector(11 downto 0);
signal mux_timestamp_S               : std_logic_vector(15 downto 0);
signal mux_superburstnumber_S        : std_logic_vector(30 downto 0);
signal mux_data_out_read_S           : std_logic;
signal mux_data_out_available_S      : std_logic;

signal pulse_channel_S               : std_logic_vector(15 downto 0);
signal pulse_statusbyte_S            : std_logic_vector(7 downto 0);
signal pulse_energy_S                : std_logic_vector(15 downto 0);
signal pulse_timefraction_S          : std_logic_vector(11 downto 0);
signal pulse_timestamp_S             : std_logic_vector(15 downto 0);
signal pulse_superburstnumber_S      : std_logic_vector(30 downto 0);

signal pulse_packet_write_S          : std_logic;
signal pulse_packet_request_S        : std_logic;
signal pulse_packet_read_S           : std_logic;
signal pulse_packet_available_S      : std_logic;
signal pulse_data_read_after1clk_S   : std_logic;

signal data64_pulse_packet_available_S : std_logic;
signal data64_wave_in_available_S    : std_logic;
signal wave_in_read_S                : std_logic;

signal combine_pulse_S               : std_logic_vector((NROFFIBERS*NROFADCS)/(2*(ADCINDEXSHIFT+1))-1 downto 0) := (others => '0');

		
signal muxstat_outfifo_fullness_S    : array_fiber16bits_type := (others => (others => '0'));
signal pulse_infifo_maxfullness_S    : array_fiber16bits_type := (others => (others => '0'));
signal muxstat_infifo_fullness_S     : array_fiber16bits_type := (others => (others => '0'));
signal pulse_outfifo_fullness_S      : std_logic_vector (15 downto 0) := (others => '0');
signal wave_infifo_fullness_S        : array_fiber16bits_type := (others => (others => '0'));
signal wave_outfifo_fullness_S       : std_logic_vector (15 downto 0) := (others => '0');
signal SelectWaveMUXfullness_S       : std_logic := '0';
signal SelectWaveMUXfullness_sync_S  : std_logic;

signal latestsuperburst_write_S      : std_logic := '0';
signal latestsuperburstnumber_S      : std_logic_vector (30 downto 0) := (others => '0');

signal timestamperrors_S             : array_fiber10bits_type := (others => (others => '0'));
signal skipped_pulses_S              : array_fiber10bits_type := (others => (others => '0'));
signal dataerrors_S                  : array_fiber10bits_type := (others => (others => '0'));
signal pulsemux_error_S              : std_logic;
signal wavemux_error_S               : std_logic;
signal pulsemux_error1_S             : std_logic;
signal wavemux_error1_S              : std_logic;
signal multiplexer_error_S           : std_logic;
signal clearerrors_S                 : std_logic_vector(0 to NROFFIBERS-1);
signal clearerrors_all_S             : std_logic;
signal clearerrors_sync_S            : std_logic;

-- SlowControl to/from cpu
signal IO_serialdata_S               : std_logic_vector(0 to NROFFIBERS-1) := (others => '0');
signal IO_serialavailable_S          : std_logic_vector(0 to NROFFIBERS-1) := (others => '0');
signal IO_byte_S                     : std_logic_vector (7 downto 0);
signal IO_write_S                    : std_logic; 

signal board_status_S                : array_muxregister_type := (others => (others => '0'));
signal board_status_read_S           : std_logic_vector(0 to NROFMUXREGS-1);
signal board_control_S               : array_muxregister_type := (others => (others => '0'));
signal board_control_write_S         : std_logic_vector(0 to NROFMUXREGS-1);

signal SODA_enable0_S                : std_logic;	

signal extractdata_start_S           : std_logic := '0';	
signal extractdata_make_selection_S  : std_logic := '0';	
signal extractdata_bothgain_S        : std_logic := '0';
signal extractdata_adcnumber_S       : std_logic_vector(15 downto 0);	
signal extractdata_ready_S           : std_logic := '0';	
signal extractdata_after1clk_ready_S : std_logic := '0';	
signal extractdata_after1clk_ready0_S : std_logic := '0';	
signal extractdata_select_S          : std_logic_vector(1 downto 0);
signal extractdata_data_S            : std_logic_vector(31 downto 0);

signal extractwave_start_S           : std_logic := '0';	
signal extractwave_make_selection_S  : std_logic := '0';	
signal extractwave_bothgain_S        : std_logic := '0';	
signal extractwave_adcnumber_S       : std_logic_vector(15 downto 0);	
signal extractwave_ready_S           : std_logic := '0';
signal extractwave_after1clk_ready_S : std_logic := '0';
signal extractwave_after1clk_ready0_S : std_logic := '0';
signal extractwave_data_read_S       : std_logic := '0';	
signal extractwave_data_S            : std_logic_vector(31 downto 0);
	
signal check_error_S                 : std_logic_vector(0 to NROFFIBERS-1);
signal wave_data_read_prev_S         : std_logic := '0';	
signal check_error2_S                : std_logic := '0';	
		
signal testword0_S                   : array_fiber36bits_type := (others => (others => '0'));
signal testword1_S                   : array_fiber36bits_type := (others => (others => '0'));
signal testword2_S                   : array_fiber36bits_type := (others => (others => '0'));
signal testPin_S                     : array_fiber4bits_type := (others => (others => '0'));

begin

process(slowcontrol_clock)
variable counter_V : integer range 0 to 7 := 0;
begin
	if (rising_edge(slowcontrol_clock)) then 
		reset_slowcontrolclock_s <= reset;
	end if;
end process;
process(packet_in_clock)
begin
	if (rising_edge(packet_in_clock)) then 
		reset_packet_in_clock_S <= reset;
	end if;
end process;
process(packet_out_clock)
begin
	if (rising_edge(packet_out_clock)) then 
		reset_packet_out_clock_S <= reset;
	end if;
end process;

		
DC_slow_control_TRB3_1: DC_slow_control_TRB3 port map(
		rst => reset_slowcontrolclock_S,
		clk => slowcontrol_clock,
		BUS_READ_IN => BUS_READ_IN,
		BUS_WRITE_IN => BUS_WRITE_IN,
		BUS_BUSY_OUT => BUS_BUSY_OUT,
		BUS_ACK_OUT => BUS_ACK_OUT,
		BUS_ADDR_IN => BUS_ADDR_IN,
		BUS_DATA_IN => BUS_DATA_IN,
		BUS_DATA_OUT => BUS_DATA_OUT,
		
		io_data_in => IO_serialdata_S,
		IO_data_in_available => IO_serialavailable_S,
		io_data_out => IO_byte_S,
		io_write_out => IO_write_S,

		extract_data_available => extractdata_after1clk_ready_S,
		extract_wave_available => extractwave_after1clk_ready_S,

		board_status => board_status_S,
		board_status_read => board_status_read_S,
		board_control => board_control_S,
		board_control_write => board_control_write_S,
		testword0 => open);

		
-- ADDRESS_MUX_FIBERMODULE_STATUS : adr=0 in MUX_fibermodule_interface
-- ADDRESS_MUX_SLOWCONTROL_SKIPPED : adr=1 not used anymore
-- ADDRESS_MUX_MULTIPLEXER_STATUS : adr=2 in MUX_fibermodule_interface

-- ADDRESS_MUX_SODA_CONTROL : adr=3 
SODA_enable0_S <= board_control_S(conv_integer(ADDRESS_MUX_SODA_CONTROL(3 downto 0)))(0);
-- not used anymore reset_timestampcounter0_S <= board_control_S(conv_integer(ADDRESS_MUX_SODA_CONTROL(3 downto 0)))(1);
EnableOutputFibre0_S <= board_control_S(conv_integer(ADDRESS_MUX_SODA_CONTROL(3 downto 0)))(4);
EnableWaveformSending_S <= board_control_S(conv_integer(ADDRESS_MUX_SODA_CONTROL(3 downto 0)))(5);
SelectWaveMUXfullness_S <= board_control_S(conv_integer(ADDRESS_MUX_SODA_CONTROL(3 downto 0)))(6);
EnableExternalSODA <= board_control_S(conv_integer(ADDRESS_MUX_SODA_CONTROL(3 downto 0)))(7);
reset_fibers0_S <= board_control_S(conv_integer(ADDRESS_MUX_SODA_CONTROL(3 downto 0)))(8);
no_packet_limit <= board_control_S(conv_integer(ADDRESS_MUX_SODA_CONTROL(3 downto 0)))(9);
DC_posedge_to_pulse_resetfibers: DC_posedge_to_pulse port map(
    clock_in => slowcontrol_clock,
    clock_out => SODA_clock,
    en_clk => '1',
    signal_in => reset_fibers0_S,
    pulse => reset_fibers);

-- ADDRESS_MUX_TIMESTAMP_ERRORS : adr=5 in MUX_fibermodule_interface


-- ADDRESS_MUX_EXTRACTWAVE : adr=7
extractwave_start_S <= board_control_write_S(conv_integer(ADDRESS_MUX_EXTRACTWAVE(3 downto 0)));
extractwave_adcnumber_S <= board_control_S(conv_integer(ADDRESS_MUX_EXTRACTWAVE(3 downto 0)))(15 downto 0);
extractwave_make_selection_S <= board_control_S(conv_integer(ADDRESS_MUX_EXTRACTWAVE(3 downto 0)))(16);
extractwave_bothgain_S <= board_control_S(conv_integer(ADDRESS_MUX_EXTRACTWAVE(3 downto 0)))(17);
board_status_S(conv_integer(ADDRESS_MUX_EXTRACTWAVE(3 downto 0))) 
	<= ones(31 downto 0) when extractwave_after1clk_ready_S='0' else extractwave_data_S;
extractwave_data_read_S <= '1' when (board_status_read_S(conv_integer(ADDRESS_MUX_EXTRACTWAVE(3 downto 0)))='1') and (extractwave_ready_S='1') else '0';

extractwave_after1clk_ready_S <= '1' when (extractwave_after1clk_ready0_S='1') and (extractwave_start_S='0') else '0';
process(slowcontrol_clock)
variable counter_V : integer range 0 to 7 := 0;
begin
	if (rising_edge(slowcontrol_clock)) then 
		if extractwave_start_S='1' then
			counter_V := 0;
			extractwave_after1clk_ready0_S <= '0';
		elsif counter_V<7 then
			counter_V := counter_V+1;
			extractwave_after1clk_ready0_S <= '0';
		else
			extractwave_after1clk_ready0_S <= extractwave_ready_S;
		end if;
	end if;
end process;

-- ADDRESS_MUX_EXTRACTDATA : adr=8
extractdata_start_S <= board_control_write_S(conv_integer(ADDRESS_MUX_EXTRACTDATA(3 downto 0)));
extractdata_adcnumber_S <= board_control_S(conv_integer(ADDRESS_MUX_EXTRACTDATA(3 downto 0)))(15 downto 0);
extractdata_make_selection_S <= board_control_S(conv_integer(ADDRESS_MUX_EXTRACTDATA(3 downto 0)))(16);
extractdata_bothgain_S <= board_control_S(conv_integer(ADDRESS_MUX_EXTRACTDATA(3 downto 0)))(17);
board_status_S(conv_integer(ADDRESS_MUX_EXTRACTDATA(3 downto 0))) 
	<= ones(31 downto 0) when extractdata_after1clk_ready_S='0' else extractdata_data_S;

extractdata_after1clk_ready_S <= '1' when (extractdata_after1clk_ready0_S='1') and (extractdata_start_S='0') else '0';
process(slowcontrol_clock)
variable counter_V : integer range 0 to 7 := 0;
begin
	if (rising_edge(slowcontrol_clock)) then 
		if extractdata_start_S='1' then
			counter_V := 0;
			extractdata_after1clk_ready0_S <= '0';
		elsif counter_V<7 then
			counter_V := counter_V+1;
			extractdata_after1clk_ready0_S <= '0';
		else
			extractdata_after1clk_ready0_S <= extractdata_ready_S;
		end if;
	end if;
end process; 

-- ADDRESS_MUX_SYSMON : adr=12 not used
board_status_S(conv_integer(ADDRESS_MUX_SYSMON(3 downto 0))) <= (others => '0');
	
-- ADDRESS_MUX_CROSSSWITCH : adr=0xd
process(slowcontrol_clock)
begin
	if (rising_edge(slowcontrol_clock)) then
		if reset_slowcontrolclock_S = '1' then 	
			for i in 0 to NROFFIBERS*NROFADCS/(ADCINDEXSHIFT+1)-1 loop
				combine_pulse_S <= (others => '0');
			end loop;
		else
			if (board_control_write_S(conv_integer(ADDRESS_MUX_CROSSSWITCH(3 downto 0)))='1') then
				--for i in 0 to 31 loop
				for i in 0 to 15 loop
					combine_pulse_S(i) <= board_control_S(conv_integer(ADDRESS_MUX_CROSSSWITCH(3 downto 0)))(i);
				end loop;
			end if;
		end if;
	end if;
end process;

-- ADDRESS_BOARDNUMBER : adr=0x2000 in MUX_fibermodule_interface

process(slowcontrol_clock)
begin
	if (rising_edge(slowcontrol_clock)) then 
		if reset_slowcontrolclock_S = '1' then 	
			extractdata_select_S <= "00";
		else
			if extractdata_start_S='1' then
				extractdata_select_S <= "00";
			elsif (board_status_read_S(conv_integer(ADDRESS_MUX_EXTRACTDATA(3 downto 0)))='1') and (extractdata_after1clk_ready_S='1') then
				extractdata_select_S <= extractdata_select_S+1;
			end if;
		end if;
	end if;
end process;

SODA_sync: process(SODA_clock) -- synchronise SODA commands
begin
	if (rising_edge(SODA_clock)) then 
		if reset_SODAclock_S = '1' then
			SODA_enable <= '1';
		else
			SODA_enable <= SODA_enable0_S;
		end if;
		reset_SODAclock_S <= reset;
	end if;
end process;

DC_fiber_module_generate: for index in 0 to NROFFIBERS-1 generate
	DC_fibermodule_interface1: DC_fibermodule_interface port map(
			slowcontrol_clock => slowcontrol_clock,
			packet_clock => packet_in_clock,
			MUX_clock => MUX_clock,
			SODA_clock => SODA_clock,
			reset => reset,
			channel => conv_std_logic_vector(index,4),
			superburst_number => superburst_number,
			superburst_update => superburst_update,
	-- SlowControl to/from cpu
			IO_byte => IO_byte_S,
			IO_write => IO_write_S,
			IO_serialdata => IO_serialdata_S(index),
			IO_serialavailable => IO_serialavailable_S(index),
	-- multiplexer status
			muxstat_infifo_fullness => muxstat_infifo_fullness_S(index),
			muxstat_outfifo_fullness => muxstat_outfifo_fullness_S(index),
			timestamp_errors => timestamperrors_S(index),
			skipped_pulses => skipped_pulses_S(index),
			dataerrors => dataerrors_S(index),
			clearerrors => clearerrors_S(index),
	-- Pulse data
			channel_out => pulse_data_array_channel_S(index),
			statusbyte_out => pulse_data_array_statusbyte_S(index),
			energy_out => pulse_data_array_energy_S(index),
			timefraction_out => pulse_data_array_timefraction_S(index),
			timestamp_out => pulse_data_array_timestamp_S(index),
			superburstnumber_out => pulse_data_array_superburstnumber_S(index),					
			pulse_data_write => pulse_data_array_write_S(index),
			pulse_data_allowed => pulse_data_array_allowed_S(index),
			pulse_data_almostfull => pulse_data_array_almostfull_S(index),
	-- Wave data
			wave_data_out => wave_data_array_S(index),
			wave_data_write => wave_data_array_write_S(index),
			wave_data_out_allowed => wave_data_array_allowed_S(index),
	-- MUX tx interface signals:
			txAsyncDataWrite => fiber_data32write(index),
			txAsyncData => fiber_data32out(index),
			txEndOfAsyncData => open,
			txAsyncFifoFull => fiber_data32fifofull(index),
			txLocked => fiber_txlocked(index),
	-- MUX rx interface signals:
			rxAsyncClk => open,
			rxAsyncDataRead => fiber_data32read(index),
			rxAsyncDataPresent => fiber_data32present(index),
			rxAsyncData => fiber_data32in(index),
			rxNotInTable => fiber_rxerror(index),
			rxLocked => fiber_rxlocked(index),
	-- Testpoints
			testword0 => open,
			testword1 => open);		
end generate;


muxstat_outfifo_fullness_generate: for index in 1 to NROFFIBERS-1 generate
	muxstat_outfifo_fullness_S(index) <= (others => '0');
	timestamperrors_S(index) <= (others => '0');
	skipped_pulses_S(index) <= (others => '0');
	dataerrors_S(index) <= (others => '0');
end generate;

--debug_slowcontrol1: if not DEBUG_SLOWCONTROL generate

sync_selectmuxfullness: process(MUX_clock)
begin
	if (rising_edge(MUX_clock)) then 
		SelectWaveMUXfullness_sync_S <= SelectWaveMUXfullness_S;
	end if;
end process;
muxstat_infifo_fullness_S <= pulse_infifo_maxfullness_S when SelectWaveMUXfullness_sync_S='0' else wave_infifo_fullness_S;
muxstat_outfifo_fullness_S(0) <= pulse_outfifo_fullness_S when SelectWaveMUXfullness_sync_S='0' else wave_outfifo_fullness_S;

DC_sorting_mux1: DC_sorting_mux port map(
		inputclock => packet_in_clock,
		MUXclock => MUX_clock,
		outputclock => packet_out_clock,
		reset => reset,
		channel_in => pulse_data_array_channel_S,
		statusbyte_in => pulse_data_array_statusbyte_S,
		energy_in => pulse_data_array_energy_S,
		timefraction_in => pulse_data_array_timefraction_S,
		timestamp_in => pulse_data_array_timestamp_S,
		superburstnumber_in => pulse_data_array_superburstnumber_S,
		data_in_write => pulse_data_array_write_S,
		data_in_allowed => pulse_data_array_allowed_S,
		data_in_almostfull => pulse_data_array_almostfull_S,
		fiber_index_out => fiber_index_S,
		channel_out => mux_channel_S,
		statusbyte_out => mux_statusbyte_S,
		energy_out => mux_energy_S,
		timefraction_out => mux_timefraction_S,
		timestamp_out => mux_timestamp_S,
		superburstnumber_out => mux_superburstnumber_S,
		data_out_read => mux_data_out_read_S,
		data_out_available => mux_data_out_available_S,
		infifo_fullness => pulse_infifo_maxfullness_S,
		outfifo_fullness => pulse_outfifo_fullness_S,
		error => pulsemux_error_S,
		testword0 => open,
		testword1 => open);

DC_combine_pulses1: DC_combine_pulses port map(
		clock => packet_out_clock,
		reset => reset_packet_out_clock_S,
		combine_pulse => combine_pulse_S,
		fiber_index_in => fiber_index_S,
		channel_in => mux_channel_S,
		statusbyte_in => mux_statusbyte_S,
		energy_in => mux_energy_S,
		timefraction_in => mux_timefraction_S,
		timestamp_in => mux_timestamp_S,
		superburstnumber_in => mux_superburstnumber_S,
		data_in_read => mux_data_out_read_S,
		data_in_available => mux_data_out_available_S,
		channel_out => pulse_channel_S,
		statusbyte_out => pulse_statusbyte_S,
		energy_out => pulse_energy_S,
		timefraction_out => pulse_timefraction_S,
		timestamp_out => pulse_timestamp_S,
		superburstnumber_out => pulse_superburstnumber_S,
		data_out_read => pulse_packet_read_S,
		data_out_available => pulse_packet_available_S
		);


		
pulse_packet_read_S <= '1' when 
		((EnableOutputFibre_S='1') and (pulse_packet_request_S='1') and (pulse_packet_available_S='1')) or  
		((EnableOutputFibre_S='0') and (pulse_packet_available_S='1')) 
	else '0';
pulse_packet_write_S <= '1' when (pulse_data_read_after1clk_S='1') else '0';
data64_pulse_packet_available_S <= pulse_packet_available_S when EnableOutputFibre_S='1' else '0';

packet_read_process: process(packet_out_clock)
begin
	if (rising_edge(packet_out_clock)) then 
		if reset_packet_out_clock_S = '1' then
			pulse_data_read_after1clk_S <= '0';
		else
			pulse_data_read_after1clk_S <= pulse_packet_read_S;
		end if;
		EnableOutputFibre_S <= EnableOutputFibre0_S;
	end if;
end process;

-- DC_wavemux1: DC_wavemux port map(
		-- inputclock => packet_in_clock,
		-- MUXclock => MUX_clock,
		-- outputclock => packet_out_clock,
		-- reset => reset,
		-- data_in => wave_data_array_S,
		-- data_in_write => wave_data_array_write_S,
		-- data_in_wave_allowed => wave_data_array_allowed_S,
		-- data_out => wave_data_S,
		-- data_out_read => wave_data_read_S,
		-- data_out_available => wave_data_available_S,
		-- infifo_fullness => wave_infifo_fullness_S,
		-- outfifo_fullness => wave_outfifo_fullness_S,
		-- testword0 => open,
		-- testword1 => open,
		-- error => wavemux_error_S);

DC_sorting_wavemux1: DC_sorting_wavemux port map(
		inputclock => packet_in_clock,
		MUXclock => MUX_clock,
		outputclock => packet_out_clock,
		reset => reset,
		data_in => wave_data_array_S,
		data_in_write => wave_data_array_write_S,
		data_in_wave_allowed => wave_data_array_allowed_S,
		data_out => wave_data_S,
		data_out_read => wave_data_read_S,
		data_out_available => wave_data_available_S,
		data_out_inpipe => open,
		infifo_fullness => wave_infifo_fullness_S,
		outfifo_fullness => wave_outfifo_fullness_S,
		error => wavemux_error_S,
		testword0 => open,
		testword1 => open);

wave_data_read_S <= '1' when 
			((EnableOutputFibre_S='1') and (EnableWaveformSending_S='1') 
				and (wave_in_read_S='1') and (wave_data_available_S='1')) 
		or  
			(((EnableOutputFibre_S='0') or (EnableWaveformSending_S='0')) 
				and ((wave_data_read0_S='1') and (wave_data_available_S='1')))
	else '0';
data64_wave_in_available_S <= wave_data_available_S 
	when (EnableOutputFibre_S='1') and (EnableWaveformSending_S='1') 
	else '0';
	
process(packet_out_clock)
begin
	if (rising_edge(packet_out_clock)) then 
		if wave_data_available_S='1' then
			wave_data_read0_S <= '1';
		else
			wave_data_read0_S <= '0';
		end if;
		wave_data_in_write_S <= wave_data_read_S;
	end if;
end process;
	

sync_superburstwrite: DC_posedge_to_pulse port map(
    clock_in => SODA_clock,
    clock_out => packet_out_clock,
    en_clk => '1',
    signal_in => superburst_update,
    pulse => latestsuperburst_write_S);
	
sync_superburstwrite_process: process(packet_out_clock)
begin
	if (rising_edge(packet_out_clock)) then 
		if latestsuperburst_write_S='1' then
			latestsuperburstnumber_S <= superburst_number;
		end if;
	end if;
end process;

DC_data_wave_to_64bit1: DC_data_wave_to_64bit port map(
		clock => packet_out_clock,
		reset => reset_packet_out_clock_S,
		latestsuperburstnumber => latestsuperburstnumber_S,
		channel => pulse_channel_S,
		statusbyte => pulse_statusbyte_S,
		energy => pulse_energy_S,
		timefraction => pulse_timefraction_S,
		timestamp => pulse_timestamp_S,
		superburstnumber => pulse_superburstnumber_S,
		data_in_available => data64_pulse_packet_available_S,
		data_in_read => pulse_packet_request_S,
		wave_in => wave_data_S,
		wave_in_available => data64_wave_in_available_S,
		wave_in_read => wave_in_read_S,
		data_out_allowed => data_out_allowed,
		data_out => data_out,
		data_out_write => data_out_write,
		data_out_first => data_out_first,
		data_out_last => data_out_last,
		error => data_out_error,
		testword0 => open,
		testword1 => open);
			
DC_posedge_to_pulse3: DC_posedge_to_pulse port map(
    clock_in => slowcontrol_clock,
    clock_out => packet_out_clock,
    en_clk => '1',
    signal_in => pulsemux_error_S,
    pulse => pulsemux_error1_S);
DC_posedge_to_pulse4: DC_posedge_to_pulse port map(
    clock_in => slowcontrol_clock,
    clock_out => packet_out_clock,
    en_clk => '1',
    signal_in => wavemux_error_S,
    pulse => wavemux_error1_S);
multiplexer_error_S <= '1' when (pulsemux_error1_S='1') or (wavemux_error1_S='1') else '0';

clearerrors_all_S <= '1' when conv_integer(unsigned(clearerrors_S))/=0 else '0';
DC_posedge_to_pulse5: DC_posedge_to_pulse port map(
    clock_in => slowcontrol_clock,
    clock_out => packet_out_clock,
    en_clk => '1',
    signal_in => clearerrors_all_S,
    pulse => clearerrors_sync_S);
	
DC_check_timestamp1: DC_check_timestamp port map(
		clock => packet_out_clock,
		reset => reset_packet_out_clock_S,
		clear => clearerrors_sync_S,
		channel => pulse_channel_S,
		statusbyte => pulse_statusbyte_S,
		energy => pulse_energy_S,
		timefraction => pulse_timefraction_S,
		timestamp => pulse_timestamp_S,
		superburstnumber => pulse_superburstnumber_S,
		pulse_data_write => pulse_packet_write_S,
		multiplexer_error => multiplexer_error_S,
		timestamp_errors => timestamperrors_S(0),
		skipped_pulses => skipped_pulses_S(0),
		dataerrors => dataerrors_S(0));
	
DC_extract_data1: DC_extract_data port map(
		write_clock => packet_out_clock,
		read_clock => slowcontrol_clock,
		reset => reset,
		start => extractdata_start_S,
		make_selection => extractdata_make_selection_S,
		dualgain => extractdata_bothgain_S,
		adcnumber => extractdata_adcnumber_S,
		channel => pulse_channel_S,
		statusbyte => pulse_statusbyte_S,
		energy => pulse_energy_S,
		timefraction => pulse_timefraction_S,
		timestamp => pulse_timestamp_S,
		superburstnumber => pulse_superburstnumber_S,
		pulse_data_write => pulse_packet_write_S,
		ready => extractdata_ready_S,
		pulse_data_select => extractdata_select_S,
		pulse_data_out => extractdata_data_S,
		testword0 => open);

DC_extract_wave1: DC_extract_wave port map(
		write_clock => packet_out_clock,
		read_clock => slowcontrol_clock,
		reset => reset,
		start => extractwave_start_S,
		make_selection => extractwave_make_selection_S,
		dualgain => extractwave_bothgain_S,
		adcnumber => extractwave_adcnumber_S,
		wave_data_in => wave_data_S,
		wave_data_in_write => wave_data_in_write_S,
		ready => extractwave_ready_S,
		wave_data_out => extractwave_data_S,
		wave_data_out_read => extractwave_data_read_S,
		testword0 => open);

DC_checkwave_all: for index in 0 to NROFFIBERS-1 generate

DC_checkwave1: DC_checkwave port map(
		clock => packet_in_clock,
		reset => reset_packet_in_clock_S,
		wave_in => wave_data_array_S(index),
		wave_in_write => wave_data_array_write_S(index),
		error => check_error_S(index));

end generate;

DC_checkwave2: DC_checkwave port map(
		clock => packet_out_clock,
		reset => reset_packet_out_clock_S,
		wave_in => wave_data_S,
		wave_in_write => wave_data_read_prev_S,
		error => check_error2_S);

-- end generate; -- DEBUG_SLOWCONTROL

process(packet_out_clock)
begin
	if (rising_edge(packet_out_clock)) then 
		wave_data_read_prev_S <= wave_data_read_S;
	end if;
end process;


testword1 <= testword1_S(0);
testword2 <= (others => '0');

		
		
end Behavioral;
